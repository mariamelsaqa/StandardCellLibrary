*** SPICE deck for cell F7_Size_1_sim{sch} from library DD2_Project
*** Created on Tue Apr 12, 2022 18:51:37
*** Last revised on Tue Apr 12, 2022 19:15:32
*** Written on Tue Apr 12, 2022 19:15:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT DD2_Project__F7_Size_1 FROM CELL F7_Size_1{sch}
.SUBCKT DD2_Project__F7_Size_1 F W X Y Z
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F X net@33 gnd nmos L=0.4U W=1.6U
Mnmos@1 net@33 Z gnd gnd nmos L=0.4U W=1.6U
Mnmos@2 F X net@36 gnd nmos L=0.4U W=1.6U
Mnmos@3 F Y net@36 gnd nmos L=0.4U W=1.6U
Mnmos@4 F Z net@36 gnd nmos L=0.4U W=1.6U
Mnmos@5 net@36 W gnd gnd nmos L=0.4U W=1.6U
Mpmos@0 net@7 X F vdd pmos L=0.4U W=22.72U
Mpmos@1 net@7 Z F vdd pmos L=0.4U W=11.36U
Mpmos@2 net@5 Y net@6 vdd pmos L=0.4U W=22.72U
Mpmos@3 net@6 Z net@7 vdd pmos L=0.4U W=22.72U
Mpmos@4 vdd X net@5 vdd pmos L=0.4U W=22.72U
Mpmos@5 vdd W net@7 vdd pmos L=0.4U W=11.36U
.ENDS DD2_Project__F7_Size_1

.global gnd vdd

*** TOP LEVEL CELL: F7_Size_1_sim{sch}
XF7_Size_@0 out X Y Z W DD2_Project__F7_Size_1

* Spice Code nodes in cell cell 'F7_Size_1_sim{sch}'
Vdd vdd 0 dc 1.8
Vin X 0 pulse 0 1.8 0.1n 400p 400p 5n 10n
Vy Y 0 dc 0
Vz Z 0 dc 1.8
Vw W 0 dc 0
.trans 0 100n
cload out 0 9fF
.measure tpdr trig v(X) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf trig v(X) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.include F:\AUC\DD2\pro1\model.txt
.END
