*** SPICE deck for cell F7_Size_2_sim{sch} from library DD2_Project
*** Created on Tue Apr 12, 2022 19:16:24
*** Last revised on Tue Apr 12, 2022 19:26:45
*** Written on Tue Apr 12, 2022 19:26:49 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT DD2_Project__F7_Size_2 FROM CELL F7_Size_2{sch}
.SUBCKT DD2_Project__F7_Size_2 F W X Y Z
** GLOBAL gnd
** GLOBAL vdd
Mnmos@6 F X net@112 gnd nmos L=0.4U W=3.2U
Mnmos@7 net@112 Z gnd gnd nmos L=0.4U W=3.2U
Mnmos@8 F X net@86 gnd nmos L=0.4U W=3.2U
Mnmos@9 F Y net@86 gnd nmos L=0.4U W=3.2U
Mnmos@10 F Z net@86 gnd nmos L=0.4U W=3.2U
Mnmos@11 net@86 W gnd gnd nmos L=0.4U W=3.2U
Mpmos@6 net@84 X F vdd pmos L=0.4U W=45.44U
Mpmos@7 net@84 Z F vdd pmos L=0.4U W=22.72U
Mpmos@8 net@129 Y net@135 vdd pmos L=0.4U W=45.44U
Mpmos@9 net@135 Z net@84 vdd pmos L=0.4U W=45.44U
Mpmos@10 vdd X net@129 vdd pmos L=0.4U W=45.44U
Mpmos@11 vdd W net@84 vdd pmos L=0.4U W=22.72U
.ENDS DD2_Project__F7_Size_2

.global gnd vdd

*** TOP LEVEL CELL: F7_Size_2_sim{sch}
XF7_Size_@0 out X Y Z W DD2_Project__F7_Size_2

* Spice Code nodes in cell cell 'F7_Size_2_sim{sch}'
Vdd vdd 0 dc 1.8
Vin X 0 pulse 0 1.8 0.1n 400p 400p 5n 10n
Vy Y 0 dc 0
Vz Z 0 dc 1.8
Vw W 0 dc 0
.trans 0 100n
cload out 0 72fF
.measure tpdr trig v(X) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf trig v(X) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.include F:\AUC\DD2\pro1\model.txt
.END
