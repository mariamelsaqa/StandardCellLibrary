*** SPICE deck for cell Inverter_Size_1_sim{sch} from library DD2_Project
*** Created on Tue Apr 12, 2022 20:09:52
*** Last revised on Tue Apr 12, 2022 20:21:38
*** Written on Tue Apr 12, 2022 20:21:41 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT DD2_Project__Inverter_Size_1 FROM CELL Inverter_Size_1{sch}
.SUBCKT DD2_Project__Inverter_Size_1 F X
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F X gnd gnd nmos L=0.4U W=0.8U
Mpmos@0 vdd X F vdd pmos L=0.4U W=5.68U
.ENDS DD2_Project__Inverter_Size_1

.global gnd vdd

*** TOP LEVEL CELL: Inverter_Size_1_sim{sch}
XInverter@0 out X DD2_Project__Inverter_Size_1

* Spice Code nodes in cell cell 'Inverter_Size_1_sim{sch}'
Vdd vdd 0 dc 1.8
Vin X 0 pulse 0 1.8 0.1n 400p 400p 5n 10n
.trans 0 100n
cload out 0 9fF
.measure tpdr trig v(X) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf trig v(X) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.include F:\AUC\DD2\pro1\model.txt
.END
